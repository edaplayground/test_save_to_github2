module M;

  initial
    $Display("M");

endmodule
